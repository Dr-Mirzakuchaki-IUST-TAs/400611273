-------------SPI-------------
-----Niloufar Dabaghi Daryan/400611273------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity SPI is
end SPI;

architecture Behavioral of SPI is

begin


end Behavioral;

